`timescale 1ps / 1ps

module simple_fpga_cvs(
    input clock
    );
endmodule

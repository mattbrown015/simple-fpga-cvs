`timescale 1ps / 1ps

module simple_fpga_cvs(
    input wire in1,
    output wire out1,
    input wire in2,
    output wire out2,
    input wire in3,
    output wire out3,
    input wire in4,
    output wire out4,
    input wire in5,
    output wire out5
    );

    assign out1 = in1;
    assign out2 = in2;
    assign out3 = in3;
    assign out4 = in4;
    assign out5 = in5;
endmodule
